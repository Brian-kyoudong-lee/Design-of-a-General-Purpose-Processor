LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY sseg IS
PORT(		bcd : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			neg : IN STD_LOGIC;
			leds, sign : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END sseg;

ARCHITECTURE Behaviour of sseg IS
	BEGIN
	PROCESS (bcd,neg)
		BEGIN
		IF neg = '0' THEN
			sign <= NOT("0000000");
		ELSE
			sign <= NOT("0000001");
		END IF;
		
		CASE bcd IS						 -- abcdefg
			WHEN "0000" => leds <= NOT("1111110");
			WHEN "0001" => leds <= NOT("0110000");
			WHEN "0010" => leds <= NOT("1101101");
			WHEN "0011" => leds <= NOT("1111001");
			WHEN "0100" => leds <= NOT("0110011");
			WHEN "0101" => leds <= NOT("1011011");
			WHEN "0110" => leds <= NOT("1011111");
			WHEN "0111" => leds <= NOT("1110000");
			WHEN "1000" => leds <= NOT("1111111");
			WHEN "1001" => leds <= NOT("1110011");
			WHEN OTHERS => leds <= NOT("0000000");
			END CASE;
		END PROCESS;
End Behaviour;